
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library axi_filter_dma_v1_00_a;
use axi_filter_dma_v1_00_a.all;


--! This component manages a BRAM storages for labeled regions.

--! The component supports different operations for creating new regions and manipulating existing ones.
--! In detail, the following operations are supported:
--!  * Create a new feature
--!  * Update an existing feature by adding an additional run
--!  * Merge two existing features
--!
--! This component is piloted by label_selection based on the runs generated by rle.
--! The results can be read out from the internal BRAM using the #FEATURE_BRAM_READOUT and #FEATURE_BRAM_RADDR ports.
--! @see label_selection
--! @see rle
entity feature_calculation is
    generic(
        ROW_LENGTH                  : positive := 640;  --! Length of a row in the input image
        ROW_LENGTH_WIDTH            : positive := 10; --! Bitwidth of #ROW_LENGTH
        NUMBER_OF_ROWS              : positive := 480;--! Number of rows in the input image
        ROW_NUMBER_WIDTH            : positive := 9;  --! Bitwidth of #NUMBER_OF_ROWS
        MAX_NUMBER_LABELS           : positive := 2045;--! Maximum number of supported labels
        FEATURE_BRAM_ADDR_WIDTH     : positive := 11  --! Address width for the BRAM holding the detected regions
    );
    port(
        clk                         : in std_logic; --! clock input
        rstn                        : in std_logic; --! negated asynchronous reset
        run_label_1                 : in std_logic_vector(FEATURE_BRAM_ADDR_WIDTH-1 downto 0);  --! Label of the region to operate on
        run_label_2                 : in std_logic_vector(FEATURE_BRAM_ADDR_WIDTH-1 downto 0);  --! A second label which is used in case of a merge operation to specify the region which shall be merged to the one with label #RUN_LABEL_1.

        start_pos                   : in std_logic_vector(ROW_LENGTH_WIDTH-1 downto 0); --! Start pos of the run which should be added to the region with #RUN_LABEL_1
        end_pos                     : in std_logic_vector(ROW_LENGTH_WIDTH-1 downto 0); --! End pos of the run which should be added to the region with #RUN_LABEL_1
        row_number                  : in std_logic_vector(ROW_NUMBER_WIDTH-1 downto 0); --! Row number of the run which should be added to the region with #RUN_LABEL_1
        update                      : in std_logic; --! set to '1' to perform an "update" operation
        merge                       : in std_logic; --! set to '1' to perform a "merge" operation
        new_feature                 : in std_logic; --! set to '1' to perform a "new feature" operation

        feature_bram_readout        : in std_logic; --! enables the feature BRAM readout. Should only be set to '1' if all image processing steps have been completed (#IDLE = '1').
        feature_bram_raddr          : in std_logic_vector(FEATURE_BRAM_ADDR_WIDTH-1 downto 0); --! Read addres for the feature BRAM
        feature_bram_left_border    : out std_logic_vector(ROW_LENGTH_WIDTH-1 downto 0); --! Left border of the feature stored at the current BRAM address #FEATURE_BRAM_RADDR
        feature_bram_right_border   : out std_logic_vector(ROW_LENGTH_WIDTH-1 downto 0); --! Right border of the feature stored at the current BRAM address #FEATURE_BRAM_RADDR
        feature_bram_upper_border   : out std_logic_vector(ROW_NUMBER_WIDTH-1 downto 0); --! Upper border of the feature stored at the current BRAM address #FEATURE_BRAM_RADDR
        feature_bram_lower_border   : out std_logic_vector(ROW_NUMBER_WIDTH-1 downto 0); --! Lower border of the feature stored at the current BRAM address #FEATURE_BRAM_RADDR
        feature_bram_valid          : out std_logic --! indicates if the feature at the current BRAM address #FEATURE_BRAM_RADDR is valid. Invalid features should be ignored.
    );
end feature_calculation;

architecture behavioral of feature_calculation is

    type FEATURE_TYPE_BOUNDS is
    record
        left, right  : std_logic_vector(ROW_LENGTH_WIDTH-1 downto 0);
        upper, lower : std_logic_vector(ROW_NUMBER_WIDTH-1 downto 0);
    end record;


    constant DATA_WIDTH_BOUNDS : positive := ROW_LENGTH_WIDTH*2 + ROW_NUMBER_WIDTH*2;

    component ram_dp is
        generic (
            ADDR_WIDTH : positive  := 2;
            DATA_WIDTH : positive  := 6;
            USE_OUTPUT_REG : std_logic  := '0'
        );
        port(
            clk : in std_logic;

            wena    : in std_logic;
            wenb    : in std_logic;
            addra   : in std_logic_vector(ADDR_WIDTH-1 downto 0);
            addrb   : in std_logic_vector(ADDR_WIDTH-1 downto 0);
            dina    : in std_logic_vector(DATA_WIDTH-1 downto 0);
            dinb    : in std_logic_vector(DATA_WIDTH-1 downto 0);
            douta   : out std_logic_vector(DATA_WIDTH-1 downto 0);
            doutb   : out std_logic_vector(DATA_WIDTH-1 downto 0)
        );
    end component;

    component ram_tp is
        generic (
            ADDR_WIDTH  : POSITIVE := 2;
            DATA_WIDTH  : POSITIVE := 6;
            USE_OUTPUT_REG : std_logic := '0'
        );
        port (
            clk             : in std_logic;
            w_addr          : in std_logic_vector(ADDR_WIDTH-1 downto 0);
            w_data          : in std_logic_vector(DATA_WIDTH-1 downto 0);
            w_enable        : in std_logic;
            r_addr_1        : in std_logic_vector(ADDR_WIDTH-1 downto 0);
            r_data_1        : out std_logic_vector(DATA_WIDTH-1 downto 0);
            r_addr_2        : in std_logic_vector(ADDR_WIDTH-1 downto 0);
            r_data_2        : out std_logic_vector(DATA_WIDTH-1 downto 0)
        );
    end component;

    signal w_enable                 : std_logic := '1';
    signal bounds_read_1            : std_logic_vector(DATA_WIDTH_BOUNDS-1 downto 0);
    signal bounds_read_2            : std_logic_vector(DATA_WIDTH_BOUNDS-1 downto 0);
    signal bounds_r_addr_1          : std_logic_vector(FEATURE_BRAM_ADDR_WIDTH-1 downto 0) := (others => '0');
    signal bounds_w_data_1          : std_logic_vector(DATA_WIDTH_BOUNDS-1 downto 0) := (others => '0');
    signal bounds_w_addr            : std_logic_vector(FEATURE_BRAM_ADDR_WIDTH-1 downto 0) := (others => '0');
    signal bounds_r_addr_2          : std_logic_vector(FEATURE_BRAM_ADDR_WIDTH-1 downto 0) := (others => '0');

    signal valid_wena               : std_logic;
    signal valid_read               : std_logic_vector(0 downto 0);
    signal valid_write              : std_logic_vector(0 downto 0);
    signal valid_read_addr          : std_logic_vector(FEATURE_BRAM_ADDR_WIDTH-1 downto 0) := (others => '0');
    signal valid_write_addr         : std_logic_vector(FEATURE_BRAM_ADDR_WIDTH-1 downto 0) := (others => '0');

-- signal bounds_1_sig, bounds_2_sig, bounds_1_before_sig, bounds_2_before_sig : FEATURE_TYPE_BOUNDS;

--READOUT Register
    signal r_readout : std_logic;

    constant max_del : integer := 2;

    type RUN_LABEL_del_type is array (natural range <>) of integer range 0 to MAX_NUMBER_LABELS;
    signal run_label_1_del, run_label_2_del :  RUN_LABEL_del_type(max_del-1 downto 0);
    signal start_pos_del, end_pos_del       :  std_logic_vector(ROW_LENGTH_WIDTH-1 downto 0);
    signal row_number_del                   : std_logic_vector(ROW_NUMBER_WIDTH-1 downto 0);
    signal update_del, merge_del, new_feature_del : std_logic_vector(max_del-1 downto 0);

begin

    bram_valid: ram_dp
    generic map(
        ADDR_WIDTH => FEATURE_BRAM_ADDR_WIDTH,
        DATA_WIDTH => 1,
        USE_OUTPUT_REG => '0'
    )
    port map(
        clk   => clk,
        addra => valid_write_addr,
        wena  => valid_wena,
        dina  => valid_write,
        douta => open,
        addrb => valid_read_addr,
        wenb  => '0',
        dinb  => (others => '0'),
        doutb => valid_read
    );


    bram_bounds: ram_tp
    generic map (
        ADDR_WIDTH => FEATURE_BRAM_ADDR_WIDTH,
        DATA_WIDTH => DATA_WIDTH_BOUNDS
    )
    port map (
        clk             => clk,
        w_addr          => bounds_w_addr,
        w_data          => bounds_w_data_1,
        w_enable        => w_enable,
        r_addr_1        => bounds_r_addr_1, --std_logiv_vector: left&right&upper&lower
        r_data_1        => bounds_read_1 ,
        r_addr_2        => bounds_r_addr_2,
        r_data_2        => bounds_read_2
    );

    bounds_r_addr_2 <= run_label_2;
    bounds_r_addr_1 <= run_label_1 when feature_bram_readout = '0' else feature_bram_raddr;
    bounds_w_addr <= std_logic_vector(to_unsigned(run_label_1_del(1), FEATURE_BRAM_ADDR_WIDTH));

    w_enable <= (merge_del(1) or update_del(1) or new_feature_del(1));

    valid_read_addr <= RUN_LABEL_1 when feature_bram_readout = '0' else feature_bram_raddr;
    valid_wena <= merge_del(1) or update_del(1) or new_feature_del(1);


    READOUT_REG : process(clk, FEATURE_BRAM_READOUT)
    begin
        if rising_edge(clk) then
            r_readout <= feature_bram_readout;
        end if;
    end process;

    UPDATE_FEATURE_SYNCHRON : process(clk, rstn, update, feature_bram_readout)
        variable addr      : integer range 0 to MAX_NUMBER_LABELS;
        variable bounds_1  : FEATURE_TYPE_BOUNDS;
        variable bounds_2  : FEATURE_TYPE_BOUNDS;

        variable valid : std_logic;
    begin

        if rstn = '0' then
            feature_bram_left_border  <= (others => '0');
            feature_bram_right_border <= (others => '0');
            feature_bram_upper_border <=(others => '0');
            feature_bram_lower_border <=(others => '0');
            feature_bram_valid <= '0';

            run_label_1_del <= (others => 0);
            run_label_2_del <= (others => 0);
            start_pos_del   <= (others => '0');
            end_pos_del     <= (others => '0');
            ROW_NUMBER_del  <= (others => '0');
            update_del      <= (others => '0');
            merge_del       <= (others => '0');
            new_feature_del <= (others => '0');

            bounds_w_data_1 <= (others => '0');

            valid := '0';
            valid_write_addr  <= (others => '0');

        elsif (rising_edge(clk)) then
            run_label_1_del(0) <= to_integer(unsigned(run_label_1));
            run_label_2_del(0) <= to_integer(unsigned(run_label_2));
            start_pos_del   <= start_pos;
            end_pos_del     <= end_pos;
            ROW_NUMBER_del  <= row_number;
            update_del(0)      <= update;
            merge_del(0)       <= merge;
            new_feature_del(0) <= new_feature;

            G0: for i in max_del-1 downto 1 loop
                run_label_1_del(i) <= run_label_1_del(i-1);
                run_label_2_del(i) <= run_label_1_del(i-1);
                update_del(i)      <= update_del(i-1);
                merge_del(i)       <= merge_del(i-1) ;
                new_feature_del(i) <= new_feature_del(i-1);
            end loop;

            bounds_w_data_1 <= (others => '0');

            if (r_readout = '1') then
                feature_bram_left_border <= bounds_read_1(DATA_WIDTH_BOUNDS-1 downto DATA_WIDTH_BOUNDS - ROW_LENGTH_WIDTH);
                feature_bram_right_border <= bounds_read_1(DATA_WIDTH_BOUNDS - ROW_LENGTH_WIDTH-1 downto DATA_WIDTH_BOUNDS - 2*ROW_LENGTH_WIDTH);
                feature_bram_upper_border <= bounds_read_1(DATA_WIDTH_BOUNDS - 2*ROW_LENGTH_WIDTH-1 downto DATA_WIDTH_BOUNDS - 2*ROW_LENGTH_WIDTH - ROW_NUMBER_WIDTH);
                feature_bram_lower_border <= bounds_read_1(DATA_WIDTH_BOUNDS - 2*ROW_LENGTH_WIDTH - ROW_NUMBER_WIDTH-1 downto 0);
                feature_bram_valid <= valid_read(0);
            end if;


            valid := valid_read(0);

            bounds_1.left  := bounds_read_1(DATA_WIDTH_BOUNDS                    - 1 downto DATA_WIDTH_BOUNDS -     ROW_LENGTH_WIDTH);
            bounds_1.right := bounds_read_1(DATA_WIDTH_BOUNDS - ROW_LENGTH_WIDTH - 1 downto DATA_WIDTH_BOUNDS - 2 * ROW_LENGTH_WIDTH);
            bounds_1.upper := bounds_read_1(DATA_WIDTH_BOUNDS - 2*ROW_LENGTH_WIDTH-1 downto DATA_WIDTH_BOUNDS - 2 * ROW_LENGTH_WIDTH - ROW_NUMBER_WIDTH);
            bounds_1.lower := bounds_read_1(DATA_WIDTH_BOUNDS - 2*ROW_LENGTH_WIDTH - ROW_NUMBER_WIDTH-1 downto 0);

            bounds_2.left  := bounds_read_2(DATA_WIDTH_BOUNDS-1                                           downto DATA_WIDTH_BOUNDS - ROW_LENGTH_WIDTH);
            bounds_2.right := bounds_read_2(DATA_WIDTH_BOUNDS-1 -   ROW_LENGTH_WIDTH                      downto DATA_WIDTH_BOUNDS - 2*ROW_LENGTH_WIDTH);
            bounds_2.upper := bounds_read_2(DATA_WIDTH_BOUNDS-1 - 2*ROW_LENGTH_WIDTH                      downto DATA_WIDTH_BOUNDS - 2*ROW_LENGTH_WIDTH - ROW_NUMBER_WIDTH);
            bounds_2.lower := bounds_read_2(DATA_WIDTH_BOUNDS   - 2*ROW_LENGTH_WIDTH - ROW_NUMBER_WIDTH-1 downto 0);

             -- bounds_1_before_sig <= bounds_1; -- useless is delayed by one clock...
             -- bounds_2_before_sig <= bounds_2;

            if update_del(0) = '1' then
                -- update left bound
                if start_pos_del < bounds_1.left then
                    bounds_1.left := start_pos_del;
                end if;
                -- update right bound
                if end_pos_del > bounds_1.right then
                    bounds_1.right := end_pos_del;
                -- set upper bound, if new label
                end if;

                if (valid ='0') then
                    bounds_1.upper := row_number_del;

                    valid := '1';

                end if;
                valid_write_addr <= std_logic_vector(to_unsigned(run_label_1_del(0), FEATURE_BRAM_ADDR_WIDTH));
                -- set lower bound, trivial
                bounds_1.lower := row_number_del;

            elsif merge_del(0) = '1' then
                -- merge left bound
                if bounds_1.left > bounds_2.left then
                    bounds_1.left := bounds_2.left;
                end if;
               -- merge right bound
                if bounds_1.right < bounds_2.right then
                    bounds_1.right := bounds_2.right;
                end if;
                -- merge upper bound
                if bounds_1.upper > bounds_2.upper then
                    bounds_1.upper := bounds_2.upper;
                end if;
               -- merge lower bound
                if bounds_1.lower < bounds_2.lower then
                    bounds_1.lower := bounds_2.lower;
                end if;

                if run_label_1_del(0) = run_label_2_del(0) then
                    valid := '1';
                else
                    valid := '0';
                end if;

                valid_write_addr <= std_logic_vector(to_unsigned(run_label_2_del(0), FEATURE_BRAM_ADDR_WIDTH));

            elsif new_feature_del(0) = '1' then
                -- set up all information of new label
                bounds_1.left :=  start_pos_del;
                bounds_1.right := end_pos_del;
                bounds_1.upper := row_number_del;
                bounds_1.lower := row_number_del;

                valid := '1';
                valid_write_addr <= std_logic_vector(to_unsigned(run_label_1_del(0), FEATURE_BRAM_ADDR_WIDTH));
            end if;

            if update_del(0) = '1' or merge_del(0) = '1' or new_feature_del(0) = '1' then
                bounds_w_data_1 <= bounds_1.left & bounds_1.right & bounds_1.upper & bounds_1.lower;
                valid_write(0) <= valid;
            end if;
        end if;

   -- bounds_1_sig <= bounds_1;
   -- bounds_2_sig <= bounds_2;

    end process;

end behavioral;

